module top_module( 
    input  logic [2:0] a, b,
    input  logic 	   cin,
    output logic [2:0] cout,
    output logic [2:0] sum );

endmodule
